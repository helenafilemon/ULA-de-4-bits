module divisor(A, B, S, Error);
    input [3:0] A, B;
    output [3:0] S;
    output Error;
    wire [3:0] nB;

    not (nB[0], B[0]);
    not (nB[1], B[1]);
    not (nB[2], B[2]);
    not (nB[3], B[3]);

    and (Error, nB[3], nB[2], nB[1], nB[0]);

  
    divisor0 (.A(A), .B(B), .S0(S[0]));
    divisor1 (.A(A), .B(B), .S1(S[1]));
    divisor2 (.A(A), .B(B), .S2(S[2]));
    divisor3 (.A(A), .B(B), .S3(S[3]));
endmodule

//=============== SUBMÓDULOS ===============

module divisor0 (A, B, S0);
    input [3:0] A, B;
    output S0;
    wire [3:0] nA, nB;
    wire [32:0] w;

    not (nA[0], A[0]);
    not (nA[1], A[1]);
    not (nA[2], A[2]);
    not (nA[3], A[3]);
    not (nB[0], B[0]);
    not (nB[1], B[1]);
    not (nB[2], B[2]);
    not (nB[3], B[3]);
            
   
    and (w[0], A[0], nB[3], nB[2], nB[1], B[0]);
    and (w[1], A[1], nB[3], nB[2], B[1], nB[0]);
    and (w[2], A[1], nA[0], nB[3], nB[2], B[1], nB[0]);
    and (w[3], nA[2], A[1], A[0], nB[3], nB[2], B[1]);
    and (w[4], nA[3], A[2], nA[1], nA[0], nB[3], nB[2], B[1], B[0]);
    and (w[5], A[2], nA[1], nB[3], B[2], nB[1], nB[0]);
    and (w[6], A[2], nA[0], nB[3], B[2], nB[1], nB[0]);
    and (w[7], nA[3], A[2], nA[1], A[0], nB[3], nB[2], B[0]);
    and (w[8], nA[3], A[2], nA[1], A[0], nB[3], B[2], nB[1]);
    and (w[9], nA[3], A[2], A[1], nA[0], nB[3], B[2], nB[1]);
    and (w[10], nA[3], A[2], A[1], nB[3], B[2], B[1], nB[0]);
    and (w[11], nA[3], A[2], A[1], A[0], nB[3], B[2]);
    and (w[12], A[2], A[1], A[0], nB[3], B[2], nB[1]);
    and (w[13], A[3], nA[2], nA[1], nB[3], B[2], B[0]);
    and (w[14], A[3], nA[2], nB[3], B[2], B[1]);
    and (w[15], A[3], nA[2], nA[1], nB[3], B[2], B[1]);
    and (w[16], A[3], nA[1], nB[3], B[2], B[1], B[0]);
    and (w[17], A[3], nA[2], nB[3], B[2], B[1], B[0]);
    and (w[18], A[3], nA[1], nA[0], nB[3], B[2], B[1], B[0]);
    and (w[19], A[3], nA[2], B[3], nB[2], nB[1], nB[0]);
    and (w[20], A[3], nA[2], nA[1], A[0], nB[3], B[1], B[0]);
    and (w[21], A[3], nA[2], A[0], B[3], nB[2], nB[1]);
    and (w[22], A[3], nA[2], A[1], nA[0], nB[3], B[1]);
    and (w[23], A[3], A[1], B[3], nB[2], nB[1]);
    and (w[24], A[3], nA[2], A[1], B[3], nB[2], nB[0]);
    and (w[25], A[3], A[1], A[0], nB[2], B[1]);
    and (w[26], A[3], A[2], nA[1], B[3], nB[2]);
    and (w[27], A[3], A[2], nA[0], B[3], nB[2]);
    and (w[28], A[3], A[2], B[3], B[2], nB[1], nB[0]);
    and (w[29], A[3], A[2], nA[1], A[0], B[3], nB[1]);
    and (w[30], A[3], A[2], A[1], nA[0], B[3], nB[1]);
    and (w[31], A[3], A[2], A[1], B[3], B[1], nB[0]);
    and (w[32], A[3], A[2], A[1], A[0], B[3], B[0]);

    
    or (S0, w[0], w[1], w[2], w[3], w[4], w[5], w[6], w[7], w[8], w[9], w[10], w[11], w[12], w[13], w[14], w[15], w[16], w[17], w[18],
         w[19], w[20], w[21], w[22], w[23], w[24], w[25], w[26], w[27], w[28], w[29], w[30], w[31], w[32]);
endmodule


module divisor1(A, B, S1);
    input [3:0] A, B;
    output S1;
    wire [3:0] nA, nB;
    wire [14:0] w;
    
    not (nA[0],A[0]); not (nA[1],A[1]); not (nA[2],A[2]); not (nA[3],A[3]);
    not (nB[0],B[0]); not (nB[1],B[1]); not (nB[2],B[2]); not (nB[3],B[3]);
    
    and (w[0],A[1],nB[3],nB[2],nB[1],B[0]);
    and (w[1],A[1],nA[0],nB[3],nB[2],nB[1],B[0]);
    and (w[2],A[2],nB[3],nB[2],B[1],nB[0]);
    and (w[3],A[2],nA[1],nB[3],nB[2],B[1],nB[0]);
    and (w[4],A[2],nA[0],nB[3],nB[2],B[1],nB[0]);
    and (w[5],nA[3],A[2],A[1],nB[3],nB[2],B[1],B[0]);
    and (w[6],A[3],nA[2],nA[1],nB[3],nB[2],B[1],B[0]);
    and (w[7],A[3],nA[2],nB[3],B[2],nB[1],nB[0]);
    and (w[8],A[3],nA[2],A[1],nB[3],nB[2],B[0]);
    and (w[9],A[3],nA[2],A[1],nA[0],nB[3],nB[2],B[0]);
    and (w[10],A[3],A[1],nB[3],B[2],nB[1],B[0]);
    and (w[11],A[3],A[2],nA[1],nB[3],B[2],nB[1]);
    and (w[12],A[3],A[2],nB[3],B[2],B[1],nB[0]);
    and (w[13],A[3],A[2],A[1],nB[3],B[2]);
    and (w[14],A[3],A[2],A[1],nA[0],nB[3],B[2]);
    
    
    or (S1,w[0],w[1],w[2],w[3],w[4],w[5],w[6],w[7],w[8],w[9],w[10],w[11],w[12],w[13],w[14]);
endmodule


module divisor2(A, B, S2);
    input [3:0] A, B;
    output S2;
    wire [3:0] nA, nB;
    wire [7:0] w;

    not (nA[0],A[0]); not (nA[1],A[1]); not (nA[2],A[2]); not (nA[3],A[3]);
    not (nB[0],B[0]); not (nB[1],B[1]); not (nB[2],B[2]); not (nB[3],B[3]);

    and (w[0],A[2],nB[3],nB[2],nB[1],B[0]);
    and (w[1],A[2],nA[1],nB[3],nB[2],nB[1],B[0]);
    and (w[2],A[2],nA[0],nB[3],nB[2],nB[1],B[0]);
    and (w[3],A[3],nB[3],nB[2],B[1],nB[0]);
    and (w[4],A[3],nA[2],nB[3],nB[2],B[1],nB[0]);
    and (w[5],A[3],nA[1],nB[3],nB[2],B[1],nB[0]);
    and (w[6],A[3],nA[0],nB[3],nB[2],B[1],nB[0]);
    and (w[7],A[3],A[2],nB[3],nB[2],B[1],B[0]);


    or (S2,w[0],w[1],w[2],w[3],w[4],w[5],w[6],w[7]);
endmodule


module divisor3(A, B, S3);
    input [3:0] A, B;
    output S3;
    wire [3:0] nA, nB;
    wire [5:0] w;

    not (nA[0],A[0]); not (nA[1],A[1]); not (nA[2],A[2]); not (nA[3],A[3]);
    not (nB[0],B[0]); not (nB[1],B[1]); not (nB[2],B[2]); not (nB[3],B[3]);

    and (w[0],A[3],nB[3],nB[2],nB[1],B[0]);
    and (w[1],A[3],nA[2],nB[3],nB[2],nB[1],B[0]);
    and (w[2],A[3],nA[1],nB[3],nB[2],nB[1],B[0]);
    and (w[3],A[3],nA[0],nB[3],nB[2],nB[1],B[0]);
    


    or (S3,w[0],w[1],w[2],w[3]);
endmodule

